library ieee;
use ieee.std_logic_1164.all;

entity tb_adder is
	generic ( wait_time : time := 10 ns;
		  N : integer := 32);
end tb_adder;

-- architecture
architecture testbench of tb_adder is

component ripple_carry_adder is
	generic (N : integer := 32);
	port (  i_X, i_Y : in std_logic_vector(N-1 downto 0);
		i_C	 : in std_logic;
		o_S	 : out std_logic_vector(N-1 downto 0);
		o_C	 : out std_logic );
end component;


-- define signals
signal s_X, s_Y, s_Sum : std_logic_vector(N-1 downto 0);
signal s_Cin, s_Cout : std_logic;

-- map signals to ports
begin
my_adder : ripple_carry_adder
port map ( i_X => s_X,
	   i_Y => s_Y,
	   i_C => s_Cin,
	   o_S => s_Sum,
	   o_C => s_Cout );


-- begin tests
test: process begin
	
	-- test 1
	s_X <= x"00000000";
	s_Y <= x"00000001";
	s_Cin <= '0';
	wait for wait_time;
	-- Expected: s_Sum = 0x0000_0001
	--	     s_C  = 0

	-- test 2
	s_X <= x"0000000A";  -- 10
	s_Y <= x"FFFFFFFF";  -- -1
	s_Cin <= '0';
	wait for wait_time;
	-- Expected: s_Sum = 9
	--	     s_C  = 1

	-- test 3
	s_X <= x"0FFFFFFF";  -- 268,435,455
	s_Y <= x"00000001";  -- 1
	s_Cin <= '0';
	wait for wait_time;
	-- Expected: s_Sum = 0x10000000
	--	     s_C  = 0

	-- test 4
	s_X <= x"000000FF";  -- 255
	s_Y <= x"00000300";  -- 768
	s_Cin <= '0';
	wait for wait_time;
	-- Expected: s_Sum = 0x000003FF
	--	     s_C  = 0

	-- test 5
	s_X <= x"FFFFFFFF";  
	s_Y <= x"00000000"; 
	s_Cin <= '1';
	wait for wait_time;
	-- Expected: s_Sum = 0
	--	     s_C  = 1

	-- test 6
	s_X <= x"FFFFFFFF";  
	s_Y <= x"FFFFFFFF"; 
	s_Cin <= '1';
	wait for wait_time;
	-- Expected: s_Sum = 0xFFFFFFFF
	--	     s_C  = 1

	-- test 7
	s_X <= x"11111111";  
	s_Y <= x"22222222"; 
	s_Cin <= '1';
	wait for wait_time;
	-- Expected: s_Sum = 0x33333334
	--	     s_C  = 0

	-- test 8
	s_X <= x"00FFEEDD";  
	s_Y <= x"00001111"; 
	s_Cin <= '1';

	wait for wait_time;
	-- Expected: s_Sum = 0x00FFFFEF
	--	     s_C  = 0

wait;
end process;

end testbench;