-- 2 to 1 Multiplexer

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity mux2t1 is
port(
	i_D0 : in std_logic;
	i_D1 : in std_logic;
	i_S : in std_logic;
	o_O : out std_logic);
end mux2t1;

architecture structural of mux2t1 is

component andg2 is
  port(i_A          : in std_logic;
       i_B          : in std_logic;
       o_F          : out std_logic);
end component;

component org2 is
  port(i_A          : in std_logic;
       i_B          : in std_logic;
       o_F          : out std_logic);
end component;

component invg is
  port(i_A          : in std_logic;
       o_F          : out std_logic);
end component;

signal s_snot, s_D1, s_D0: std_logic;

begin
	not_s: invg port map (i_A => i_S,
				o_F => s_snot) ;

	and0: andg2 port map (i_A => i_D0,
				i_B => s_snot,
				o_F => s_D0);

	and1: andg2 port map (i_A => i_D1,
				i_B => i_S,
				o_F => s_D1);

	or_out: org2 port map (i_A => s_D0,
				i_B => s_D1,
				o_F => o_O);

end structural;
