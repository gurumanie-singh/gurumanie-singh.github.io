library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_textio.all;  -- For logic types I/O
library std;
use std.env.all;                -- For hierarchical/external signals
use std.textio.all;             -- For basic I/O

entity tb_mux2t1_N is
	generic(wait_time: time := 10 ns;
		  N: integer := 32);

end tb_mux2t1_N;

architecture mixed of tb_mux2t1_N is

component mux_32t1_n is
	generic (N : integer:= 32);
	port ( 
		i_D0, i_D1, i_D2, i_D3, i_D4, i_D5, i_D6,
		i_D7, i_D8, i_D9, i_D10, i_D11, i_D12, i_D13, i_D14, i_D15,
		i_D16, i_D17, i_D18, i_D19, i_D20, i_D21, i_D22, i_D23,
		i_D24, i_D25, i_D26, i_D27, i_D28, i_D29, i_D30, i_D31		: in std_logic_vector(N-1 downto 0);
		
		i_S : in std_logic_vector(4 downto 0);
		o_out : out std_logic_vector(N-1 downto 0));
end component;

-- define input/output signals, pre-set to 0
signal	s_D0,
	s_D1, 
	s_D2, 
	s_D3, 
	s_D4, 
	s_D5, 
	s_D6, 
	s_D7, 
	s_D8, 
	s_D9, 
	s_D10, 
	s_D11, 
	s_D12, 
	s_D13, 
	s_D14, 
	s_D15, 
	s_D16, 
	s_D17, 
	s_D18, 
	s_D19, 
	s_D20, 
	s_D21, 
	s_D22, 
	s_D23, 
	s_D24, 
	s_D25, 
	s_D26, 
	s_D27,	 
	s_D28, 
	s_D29, 
	s_D30, 
	s_D31 : std_logic_vector(N-1 downto 0);
signal s_iS: std_logic_vector(4 downto 0);
signal s_out: std_logic_vector(N-1 downto 0);

begin

-- map signals to mux ports
my_mux: mux_32t1_N
port map ( i_D0 => s_D0,
           i_D1 => s_D1,
           i_D2 => s_D2,
           i_D3 => s_D3,
           i_D4 => s_D4,
           i_D5 => s_D5,
           i_D6 => s_D6,
           i_D7 => s_D7,
           i_D8 => s_D8,
           i_D9 => s_D9,
           i_D10 => s_D10,
           i_D11 => s_D11,
           i_D12 => s_D12,
           i_D13 => s_D13,
           i_D14 => s_D14,
           i_D15 => s_D15,
           i_D16 => s_D16,
           i_D17 => s_D17,
           i_D18 => s_D18,
           i_D19 => s_D19,
           i_D20 => s_D20,
           i_D21 => s_D21,
           i_D22 => s_D22,
           i_D23 => s_D23,
           i_D24 => s_D24,
           i_D25 => s_D25,
           i_D26 => s_D26,
           i_D27 => s_D27,
           i_D28 => s_D28,
           i_D29 => s_D29,
           i_D30 => s_D30,
           i_D31 => s_D31,
	   i_S => s_iS,
	   o_out => s_out);

-- begin test cases
TEST: process
begin

-- set the values of each input
s_D0 <= x"00000000";
s_D1 <= x"00000001";
s_D2 <= x"00000002";
s_D3 <= x"00000003";
s_D4 <= x"00000004";
s_D5 <= x"00000005";
s_D6 <= x"00000006";
s_D7 <= x"00000007";
s_D8 <= x"00000008";
s_D9 <= x"00000009";
s_D10 <= x"0000000A";
s_D11 <= x"0000000B";
s_D12 <= x"0000000C";
s_D13 <= x"0000000D";
s_D14 <= x"0000000E";
s_D15 <= x"0000000F";
s_D16 <= x"00000010";
s_D17 <= x"00000011";
s_D18 <= x"00000012";
s_D19 <= x"00000013";
s_D20 <= x"00000014";
s_D21 <= x"00000015";
s_D22 <= x"00000016";
s_D23 <= x"00000017";
s_D24 <= x"00000018";
s_D25 <= x"00000019";
s_D26 <= x"0000001A";
s_D27 <= x"0000001B";
s_D28 <= x"0000001C";
s_D29 <= x"0000001D";
s_D30 <= x"0000001E";
s_D31 <= x"0000001F";

-- test each select line
s_iS <= "00000";
wait for 10 ns;

s_iS <= "00001";
wait for 10 ns;

s_iS <= "00010";
wait for 10 ns;

s_iS <= "00011";
wait for 10 ns;

s_iS <= "00100";
wait for 10 ns;

s_iS <= "00101";
wait for 10 ns;

s_iS <= "00110";
wait for 10 ns;

s_iS <= "00111";
wait for 10 ns;

s_iS <= "01000";
wait for 10 ns;

s_iS <= "01001";
wait for 10 ns;

s_iS <= "01010";
wait for 10 ns;

s_iS <= "01011";
wait for 10 ns;

s_iS <= "01100";
wait for 10 ns;

s_iS <= "01101";
wait for 10 ns;

s_iS <= "01110";
wait for 10 ns;

s_iS <= "01111";
wait for 10 ns;

s_iS <= "10000";
wait for 10 ns;

s_iS <= "10001";
wait for 10 ns;

s_iS <= "10010";
wait for 10 ns;

s_iS <= "10011";
wait for 10 ns;

s_iS <= "10100";
wait for 10 ns;

s_iS <= "10101";
wait for 10 ns;

s_iS <= "10110";
wait for 10 ns;

s_iS <= "10111";
wait for 10 ns;

s_iS <= "11000";
wait for 10 ns;

s_iS <= "11001";
wait for 10 ns;

s_iS <= "11010";
wait for 10 ns;

s_iS <= "11011";
wait for 10 ns;

s_iS <= "11100";
wait for 10 ns;

s_iS <= "11101";
wait for 10 ns;

s_iS <= "11110";
wait for 10 ns;

s_iS <= "11111";
wait for 10 ns;
	
end process;

end mixed;