library IEEE;
use IEEE.std_logic_1164.all;

-- entity
entity tb_onescomp is 
	generic ( N: integer := 32;
		  wait_time: time := 10 ns);
end tb_onescomp;

-- architecture
architecture structural of tb_onescomp is

-- onescomp component
component onescomp is
	generic ( N: integer := 32);
	port ( i_in: in std_logic_vector(N-1 downto 0);
	       o_O: out std_logic_vector(N-1 downto 0));
end component;

-- define signals
signal s_in, s_out: std_logic_vector(N-1 downto 0);

-- link signals to ports
begin
my_onescomp: onescomp
port map ( i_in => s_in,
	   o_O => s_out);


-- start tests
tests: process begin

-- test 1
s_in <= x"FFFFFFFF";
wait for wait_time;
-- Expected: s_out = 0x0000_0000

-- test 2
s_in <= x"00000001";
wait for wait_time;
-- Expected: s_out = 0xFFFF_FFFE

-- test 3
s_in <= x"000F000F";
wait for wait_time;
-- Expected: s_out = 0xFFF0_FFF0

-- test 4
s_in <= x"FEDCBA98";
wait for wait_time;
-- Expected: s_out = 0x0123_4567

-- test 5
s_in <= x"76543210";
wait for wait_time;
-- Expected: s_out = 0x89AB_CDEF

-- test 6
s_in <= x"05310FF2";
wait for wait_time;
-- Expected: s_out = 0xFACE_F00D

end process;

end structural;

	